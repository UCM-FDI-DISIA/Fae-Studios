sanctuaryID 0
lifeShards 0 _
earth 1
water 1
fire 1
map_key earthMap 0
earth_boss 0
water_boss 0
fire_boss 0
earth_map_rooms 0 1 1 1 2 1 3 0 4 1 5 1 6 1 7 0 8 0 9 0 10 0 11 0 12 0 13 1 14 0 15 0 16 0 17 0 18 0 19 0 _
water_map_rooms 0 1 1 1 2 1 3 1 4 1 5 1 6 0 7 1 8 1 9 0 10 0 11 0 12 1 13 0 14 0 15 0 16 0 17 0 18 0 19 0 _
fire_map_rooms 0 1 1 0 2 0 3 0 4 0 5 0 6 0 7 0 8 0 9 0 10 0 11 0 12 0 13 0 14 0 15 0 16 0 17 0 18 0 19 0 _
