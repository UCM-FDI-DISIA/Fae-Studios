sanctuaryID 0
lifeShards 1 3 _
earth 1
water 1
fire 1
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 0 2 0 3 0 4 0 5 0 6 0 7 0 8 0 9 0 10 0 11 0 12 0 13 0 14 1 15 1 16 0 17 1 18 1 19 1 20 1 21 1 22 1 23 1 24 0 25 0 26 1 27 0 _
water_map_rooms _
fire_map_rooms _
