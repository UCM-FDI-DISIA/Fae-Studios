sanctuaryID 0
lifeShards 1 3 _
earth 1
water 1
fire 1
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 0 2 0 3 0 4 0 5 0 6 0 7 0 8 0 9 0 10 0 11 0 12 0 13 0 14 1 15 0 16 0 17 0 18 0 19 0 20 0 21 0 22 0 23 0 24 0 25 0 26 0 27 0 28 1 29 1 30 0 31 1 32 1 33 1 34 1 35 1 36 1 37 1 38 0 39 0 40 1 41 0 _
water_map_rooms _
fire_map_rooms _
