sanctuaryID 0
lifeShards 0 _
earth 1
water 0
fire 0
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 1 2 1 3 0 4 0 5 0 6 1 7 1 8 0 9 0 10 0 11 0 12 0 13 0 _
water_map_rooms 0 1 1 0 2 0 3 0 4 0 5 0 6 0 7 0 8 0 9 0 10 0 11 0 12 0 _
fire_map_rooms _
