sanctuaryID 3
lifeShards 1 1 _
earth 1
water 1
fire 1
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 1 2 1 3 1 4 1 5 0 6 1 7 0 8 0 9 0 10 0 11 0 12 1 13 1 14 1 15 0 16 0 17 0 18 0 19 0 20 0 21 1 22 1 23 0 24 0 25 0 26 1 27 0 28 1 29 1 30 0 31 0 32 0 33 0 34 1 35 1 36 1 37 0 38 0 39 0 40 1 41 0 42 1 43 0 44 0 45 0 46 0 47 0 48 0 49 1 50 1 51 0 52 0 53 0 54 1 55 0 56 1 57 1 58 0 59 0 60 0 61 0 62 0 63 0 64 0 65 0 66 0 67 0 68 0 69 0 _
water_map_rooms _
fire_map_rooms _
