sanctuaryID 0
lifeShards 2 0 1 _
earth 1
water 0
fire 1
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 1 2 0 3 0 4 0 5 0 6 0 _
water_map_rooms _
fire_map_rooms _
