sanctuaryID 0
lifeShards 1 1 _
earth 1
water 1
fire 1
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 1 2 0 3 0 4 0 5 0 6 1 7 0 8 0 9 0 10 0 11 0 12 0 13 0 14 1 15 1 16 0 17 0 18 0 19 0 20 0 21 1 22 1 23 0 24 0 25 0 26 1 27 0 28 1 29 0 30 0 31 0 32 0 33 0 34 0 35 0 36 0 37 0 38 0 39 0 40 0 41 0 42 1 43 1 44 0 45 0 46 0 47 0 48 1 49 1 50 1 51 1 52 0 53 1 54 1 55 1 _
water_map_rooms _
fire_map_rooms _
