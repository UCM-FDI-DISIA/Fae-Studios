sanctuaryID 2
lifeShards 0 _
earth 1
water 1
fire 1
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 0 2 0 3 0 4 0 5 0 6 0 7 1 8 1 9 0 10 0 11 0 12 1 13 0 14 1 15 1 16 0 17 0 18 0 19 0 20 1 21 1 22 1 23 0 24 0 25 0 26 1 27 0 28 1 29 0 30 0 31 0 32 0 33 0 34 0 35 1 36 1 37 0 38 0 39 0 40 1 41 0 42 1 43 1 44 0 45 0 46 0 47 0 48 0 49 0 50 0 51 0 52 0 53 0 54 0 55 0 _
water_map_rooms _
fire_map_rooms _
