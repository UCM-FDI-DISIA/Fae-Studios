sanctuaryID 8
lifeShards 0 _
earth 1
water 1
fire 1
map_key fireMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 0 2 0 3 0 4 0 5 0 6 0 7 0 8 0 9 0 10 1 11 0 _
water_map_rooms _
fire_map_rooms _
