sanctuaryID 2
lifeShards 1 1 _
earth 1
water 1
fire 1
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 1 2 0 3 0 4 0 5 0 6 0 7 1 8 1 9 0 10 0 11 0 12 1 13 0 14 1 15 0 16 0 17 0 18 0 19 0 20 0 21 0 22 0 23 0 24 0 25 0 26 0 27 0 28 1 29 1 30 0 31 0 32 0 33 0 34 1 35 1 36 1 37 1 38 0 39 1 40 1 41 1 _
water_map_rooms _
fire_map_rooms _
