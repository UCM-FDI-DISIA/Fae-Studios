sanctuaryID 3
lifeShards 1 3 _
earth 1
water 0
fire 0
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 1 2 1 3 1 4 1 5 0 6 1 7 1 8 1 9 1 10 0 11 1 12 1 13 1 _
water_map_rooms _
fire_map_rooms _
