sanctuaryID 7
lifeShards 0 _
earth 1
water 1
fire 1
map_key waterMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 1 2 1 3 1 4 1 5 1 6 0 7 1 8 1 9 0 10 0 11 0 12 1 13 0 14 0 15 0 _
water_map_rooms _
fire_map_rooms _
