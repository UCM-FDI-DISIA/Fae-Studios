sanctuaryID 3
lifeShards 0 _
earth 1
water 1
fire 1
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 0
earth_map_rooms 0 1 1 1 2 1 3 0 4 1 5 1 6 1 7 1 8 1 9 0 10 1 11 1 12 1 13 1 _
water_map_rooms _
fire_map_rooms _
