sanctuaryID 0
lifeShards 1 3 _
earth 1
water 1
fire 1
map_key earthMap 0
earth_boss 1
water_boss 1
fire_boss 1
earth_map_rooms 0 1 1 1 2 0 3 1 4 1 5 1 6 1 7 1 8 1 9 1 10 0 11 0 12 1 13 0 14 1 15 1 16 0 17 0 18 0 19 0 20 0 21 0 22 0 23 0 24 0 25 0 26 0 27 0 _
water_map_rooms _
fire_map_rooms _
